// SoC2.v

// Generated using ACDS version 13.0 156 at 2024.10.30.12:11:00

`timescale 1 ps / 1 ps
module SoC2 (
		input  wire  clk_clk,            //         clk.clk
		input  wire  reset_reset_n,      //       reset.reset_n
		input  wire  receive_req_export, // receive_req.export
		output wire  req_export,         //         req.export
		input  wire  receive_ack_export, // receive_ack.export
		output wire  ack_export          //         ack.export
	);

	wire         nios_instruction_master_waitrequest;                                                         // NIOS_instruction_master_translator:av_waitrequest -> NIOS:i_waitrequest
	wire  [17:0] nios_instruction_master_address;                                                             // NIOS:i_address -> NIOS_instruction_master_translator:av_address
	wire         nios_instruction_master_read;                                                                // NIOS:i_read -> NIOS_instruction_master_translator:av_read
	wire  [31:0] nios_instruction_master_readdata;                                                            // NIOS_instruction_master_translator:av_readdata -> NIOS:i_readdata
	wire         nios_data_master_waitrequest;                                                                // NIOS_data_master_translator:av_waitrequest -> NIOS:d_waitrequest
	wire  [31:0] nios_data_master_writedata;                                                                  // NIOS:d_writedata -> NIOS_data_master_translator:av_writedata
	wire  [17:0] nios_data_master_address;                                                                    // NIOS:d_address -> NIOS_data_master_translator:av_address
	wire         nios_data_master_write;                                                                      // NIOS:d_write -> NIOS_data_master_translator:av_write
	wire         nios_data_master_read;                                                                       // NIOS:d_read -> NIOS_data_master_translator:av_read
	wire  [31:0] nios_data_master_readdata;                                                                   // NIOS_data_master_translator:av_readdata -> NIOS:d_readdata
	wire         nios_data_master_debugaccess;                                                                // NIOS:jtag_debug_module_debugaccess_to_roms -> NIOS_data_master_translator:av_debugaccess
	wire   [3:0] nios_data_master_byteenable;                                                                 // NIOS:d_byteenable -> NIOS_data_master_translator:av_byteenable
	wire         nios_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                           // NIOS:jtag_debug_module_waitrequest -> NIOS_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // NIOS_jtag_debug_module_translator:av_writedata -> NIOS:jtag_debug_module_writedata
	wire   [8:0] nios_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // NIOS_jtag_debug_module_translator:av_address -> NIOS:jtag_debug_module_address
	wire         nios_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // NIOS_jtag_debug_module_translator:av_write -> NIOS:jtag_debug_module_write
	wire         nios_jtag_debug_module_translator_avalon_anti_slave_0_read;                                  // NIOS_jtag_debug_module_translator:av_read -> NIOS:jtag_debug_module_read
	wire  [31:0] nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // NIOS:jtag_debug_module_readdata -> NIOS_jtag_debug_module_translator:av_readdata
	wire         nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // NIOS_jtag_debug_module_translator:av_debugaccess -> NIOS:jtag_debug_module_debugaccess
	wire   [3:0] nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // NIOS_jtag_debug_module_translator:av_byteenable -> NIOS:jtag_debug_module_byteenable
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_writedata;                                             // RAM_s1_translator:av_writedata -> RAM:writedata
	wire  [13:0] ram_s1_translator_avalon_anti_slave_0_address;                                               // RAM_s1_translator:av_address -> RAM:address
	wire         ram_s1_translator_avalon_anti_slave_0_chipselect;                                            // RAM_s1_translator:av_chipselect -> RAM:chipselect
	wire         ram_s1_translator_avalon_anti_slave_0_clken;                                                 // RAM_s1_translator:av_clken -> RAM:clken
	wire         ram_s1_translator_avalon_anti_slave_0_write;                                                 // RAM_s1_translator:av_write -> RAM:write
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_readdata;                                              // RAM:readdata -> RAM_s1_translator:av_readdata
	wire   [3:0] ram_s1_translator_avalon_anti_slave_0_byteenable;                                            // RAM_s1_translator:av_byteenable -> RAM:byteenable
	wire         jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // JTAG:av_waitrequest -> JTAG_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // JTAG_avalon_jtag_slave_translator:av_writedata -> JTAG:av_writedata
	wire   [0:0] jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // JTAG_avalon_jtag_slave_translator:av_address -> JTAG:av_address
	wire         jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // JTAG_avalon_jtag_slave_translator:av_chipselect -> JTAG:av_chipselect
	wire         jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // JTAG_avalon_jtag_slave_translator:av_write -> JTAG:av_write_n
	wire         jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // JTAG_avalon_jtag_slave_translator:av_read -> JTAG:av_read_n
	wire  [31:0] jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // JTAG:av_readdata -> JTAG_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] pcu_control_slave_translator_avalon_anti_slave_0_writedata;                                  // PCU_control_slave_translator:av_writedata -> PCU:writedata
	wire   [3:0] pcu_control_slave_translator_avalon_anti_slave_0_address;                                    // PCU_control_slave_translator:av_address -> PCU:address
	wire         pcu_control_slave_translator_avalon_anti_slave_0_write;                                      // PCU_control_slave_translator:av_write -> PCU:write
	wire  [31:0] pcu_control_slave_translator_avalon_anti_slave_0_readdata;                                   // PCU:readdata -> PCU_control_slave_translator:av_readdata
	wire         pcu_control_slave_translator_avalon_anti_slave_0_begintransfer;                              // PCU_control_slave_translator:av_begintransfer -> PCU:begintransfer
	wire   [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                  // SYSID_control_slave_translator:av_address -> SYSID:address
	wire  [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                 // SYSID:readdata -> SYSID_control_slave_translator:av_readdata
	wire   [1:0] receive_req_s1_translator_avalon_anti_slave_0_address;                                       // RECEIVE_REQ_s1_translator:av_address -> RECEIVE_REQ:address
	wire  [31:0] receive_req_s1_translator_avalon_anti_slave_0_readdata;                                      // RECEIVE_REQ:readdata -> RECEIVE_REQ_s1_translator:av_readdata
	wire   [1:0] receive_ack_s1_translator_avalon_anti_slave_0_address;                                       // RECEIVE_ACK_s1_translator:av_address -> RECEIVE_ACK:address
	wire  [31:0] receive_ack_s1_translator_avalon_anti_slave_0_readdata;                                      // RECEIVE_ACK:readdata -> RECEIVE_ACK_s1_translator:av_readdata
	wire  [31:0] req_s1_translator_avalon_anti_slave_0_writedata;                                             // REQ_s1_translator:av_writedata -> REQ:writedata
	wire   [1:0] req_s1_translator_avalon_anti_slave_0_address;                                               // REQ_s1_translator:av_address -> REQ:address
	wire         req_s1_translator_avalon_anti_slave_0_chipselect;                                            // REQ_s1_translator:av_chipselect -> REQ:chipselect
	wire         req_s1_translator_avalon_anti_slave_0_write;                                                 // REQ_s1_translator:av_write -> REQ:write_n
	wire  [31:0] req_s1_translator_avalon_anti_slave_0_readdata;                                              // REQ:readdata -> REQ_s1_translator:av_readdata
	wire  [31:0] ack_s1_translator_avalon_anti_slave_0_writedata;                                             // ACK_s1_translator:av_writedata -> ACK:writedata
	wire   [1:0] ack_s1_translator_avalon_anti_slave_0_address;                                               // ACK_s1_translator:av_address -> ACK:address
	wire         ack_s1_translator_avalon_anti_slave_0_chipselect;                                            // ACK_s1_translator:av_chipselect -> ACK:chipselect
	wire         ack_s1_translator_avalon_anti_slave_0_write;                                                 // ACK_s1_translator:av_write -> ACK:write_n
	wire  [31:0] ack_s1_translator_avalon_anti_slave_0_readdata;                                              // ACK:readdata -> ACK_s1_translator:av_readdata
	wire         nios_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios_instruction_master_translator_avalon_universal_master_0_burstcount;                     // NIOS_instruction_master_translator:uav_burstcount -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios_instruction_master_translator_avalon_universal_master_0_writedata;                      // NIOS_instruction_master_translator:uav_writedata -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] nios_instruction_master_translator_avalon_universal_master_0_address;                        // NIOS_instruction_master_translator:uav_address -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios_instruction_master_translator_avalon_universal_master_0_lock;                           // NIOS_instruction_master_translator:uav_lock -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios_instruction_master_translator_avalon_universal_master_0_write;                          // NIOS_instruction_master_translator:uav_write -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios_instruction_master_translator_avalon_universal_master_0_read;                           // NIOS_instruction_master_translator:uav_read -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios_instruction_master_translator_avalon_universal_master_0_readdata;                       // NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS_instruction_master_translator:uav_readdata
	wire         nios_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // NIOS_instruction_master_translator:uav_debugaccess -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios_instruction_master_translator_avalon_universal_master_0_byteenable;                     // NIOS_instruction_master_translator:uav_byteenable -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // NIOS_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS_instruction_master_translator:uav_readdatavalid
	wire         nios_data_master_translator_avalon_universal_master_0_waitrequest;                           // NIOS_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS_data_master_translator:uav_waitrequest
	wire   [2:0] nios_data_master_translator_avalon_universal_master_0_burstcount;                            // NIOS_data_master_translator:uav_burstcount -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios_data_master_translator_avalon_universal_master_0_writedata;                             // NIOS_data_master_translator:uav_writedata -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] nios_data_master_translator_avalon_universal_master_0_address;                               // NIOS_data_master_translator:uav_address -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios_data_master_translator_avalon_universal_master_0_lock;                                  // NIOS_data_master_translator:uav_lock -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios_data_master_translator_avalon_universal_master_0_write;                                 // NIOS_data_master_translator:uav_write -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios_data_master_translator_avalon_universal_master_0_read;                                  // NIOS_data_master_translator:uav_read -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios_data_master_translator_avalon_universal_master_0_readdata;                              // NIOS_data_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS_data_master_translator:uav_readdata
	wire         nios_data_master_translator_avalon_universal_master_0_debugaccess;                           // NIOS_data_master_translator:uav_debugaccess -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios_data_master_translator_avalon_universal_master_0_byteenable;                            // NIOS_data_master_translator:uav_byteenable -> NIOS_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios_data_master_translator_avalon_universal_master_0_readdatavalid;                         // NIOS_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS_data_master_translator:uav_readdatavalid
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // NIOS_jtag_debug_module_translator:uav_waitrequest -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> NIOS_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> NIOS_jtag_debug_module_translator:uav_writedata
	wire  [17:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> NIOS_jtag_debug_module_translator:uav_address
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> NIOS_jtag_debug_module_translator:uav_write
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> NIOS_jtag_debug_module_translator:uav_lock
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> NIOS_jtag_debug_module_translator:uav_read
	wire  [31:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // NIOS_jtag_debug_module_translator:uav_readdata -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // NIOS_jtag_debug_module_translator:uav_readdatavalid -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NIOS_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> NIOS_jtag_debug_module_translator:uav_byteenable
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // RAM_s1_translator:uav_waitrequest -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RAM_s1_translator:uav_burstcount
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RAM_s1_translator:uav_writedata
	wire  [17:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> RAM_s1_translator:uav_address
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> RAM_s1_translator:uav_write
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RAM_s1_translator:uav_lock
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> RAM_s1_translator:uav_read
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // RAM_s1_translator:uav_readdata -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // RAM_s1_translator:uav_readdatavalid -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RAM_s1_translator:uav_debugaccess
	wire   [3:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RAM_s1_translator:uav_byteenable
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // JTAG_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_avalon_jtag_slave_translator:uav_writedata
	wire  [17:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_avalon_jtag_slave_translator:uav_address
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_avalon_jtag_slave_translator:uav_write
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_avalon_jtag_slave_translator:uav_lock
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // JTAG_avalon_jtag_slave_translator:uav_readdata -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // JTAG_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // PCU_control_slave_translator:uav_waitrequest -> PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PCU_control_slave_translator:uav_burstcount
	wire  [31:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PCU_control_slave_translator:uav_writedata
	wire  [17:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> PCU_control_slave_translator:uav_address
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> PCU_control_slave_translator:uav_write
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PCU_control_slave_translator:uav_lock
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> PCU_control_slave_translator:uav_read
	wire  [31:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // PCU_control_slave_translator:uav_readdata -> PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // PCU_control_slave_translator:uav_readdatavalid -> PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PCU_control_slave_translator:uav_debugaccess
	wire   [3:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // PCU_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PCU_control_slave_translator:uav_byteenable
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // PCU_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // PCU_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // PCU_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // PCU_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // SYSID_control_slave_translator:uav_waitrequest -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SYSID_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SYSID_control_slave_translator:uav_writedata
	wire  [17:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> SYSID_control_slave_translator:uav_address
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> SYSID_control_slave_translator:uav_write
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SYSID_control_slave_translator:uav_lock
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> SYSID_control_slave_translator:uav_read
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // SYSID_control_slave_translator:uav_readdata -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // SYSID_control_slave_translator:uav_readdatavalid -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SYSID_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // SYSID_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SYSID_control_slave_translator:uav_byteenable
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // RECEIVE_REQ_s1_translator:uav_waitrequest -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] receive_req_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RECEIVE_REQ_s1_translator:uav_burstcount
	wire  [31:0] receive_req_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RECEIVE_REQ_s1_translator:uav_writedata
	wire  [17:0] receive_req_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_address -> RECEIVE_REQ_s1_translator:uav_address
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_write -> RECEIVE_REQ_s1_translator:uav_write
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RECEIVE_REQ_s1_translator:uav_lock
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_read -> RECEIVE_REQ_s1_translator:uav_read
	wire  [31:0] receive_req_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // RECEIVE_REQ_s1_translator:uav_readdata -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // RECEIVE_REQ_s1_translator:uav_readdatavalid -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RECEIVE_REQ_s1_translator:uav_debugaccess
	wire   [3:0] receive_req_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RECEIVE_REQ_s1_translator:uav_byteenable
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // RECEIVE_ACK_s1_translator:uav_waitrequest -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RECEIVE_ACK_s1_translator:uav_burstcount
	wire  [31:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RECEIVE_ACK_s1_translator:uav_writedata
	wire  [17:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_address -> RECEIVE_ACK_s1_translator:uav_address
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_write -> RECEIVE_ACK_s1_translator:uav_write
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RECEIVE_ACK_s1_translator:uav_lock
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_read -> RECEIVE_ACK_s1_translator:uav_read
	wire  [31:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // RECEIVE_ACK_s1_translator:uav_readdata -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // RECEIVE_ACK_s1_translator:uav_readdatavalid -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RECEIVE_ACK_s1_translator:uav_debugaccess
	wire   [3:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RECEIVE_ACK_s1_translator:uav_byteenable
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         req_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // REQ_s1_translator:uav_waitrequest -> REQ_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] req_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // REQ_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> REQ_s1_translator:uav_burstcount
	wire  [31:0] req_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // REQ_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> REQ_s1_translator:uav_writedata
	wire  [17:0] req_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // REQ_s1_translator_avalon_universal_slave_0_agent:m0_address -> REQ_s1_translator:uav_address
	wire         req_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // REQ_s1_translator_avalon_universal_slave_0_agent:m0_write -> REQ_s1_translator:uav_write
	wire         req_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // REQ_s1_translator_avalon_universal_slave_0_agent:m0_lock -> REQ_s1_translator:uav_lock
	wire         req_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // REQ_s1_translator_avalon_universal_slave_0_agent:m0_read -> REQ_s1_translator:uav_read
	wire  [31:0] req_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // REQ_s1_translator:uav_readdata -> REQ_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         req_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // REQ_s1_translator:uav_readdatavalid -> REQ_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         req_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // REQ_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> REQ_s1_translator:uav_debugaccess
	wire   [3:0] req_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // REQ_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> REQ_s1_translator:uav_byteenable
	wire         req_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         req_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         req_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] req_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         req_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> REQ_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // REQ_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> REQ_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // ACK_s1_translator:uav_waitrequest -> ACK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // ACK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ACK_s1_translator:uav_burstcount
	wire  [31:0] ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // ACK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ACK_s1_translator:uav_writedata
	wire  [17:0] ack_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // ACK_s1_translator_avalon_universal_slave_0_agent:m0_address -> ACK_s1_translator:uav_address
	wire         ack_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // ACK_s1_translator_avalon_universal_slave_0_agent:m0_write -> ACK_s1_translator:uav_write
	wire         ack_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // ACK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ACK_s1_translator:uav_lock
	wire         ack_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // ACK_s1_translator_avalon_universal_slave_0_agent:m0_read -> ACK_s1_translator:uav_read
	wire  [31:0] ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // ACK_s1_translator:uav_readdata -> ACK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // ACK_s1_translator:uav_readdatavalid -> ACK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // ACK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ACK_s1_translator:uav_debugaccess
	wire   [3:0] ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // ACK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ACK_s1_translator:uav_byteenable
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ACK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // ACK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ACK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // NIOS_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // NIOS_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // NIOS_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [92:0] nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // NIOS_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // NIOS_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // NIOS_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // NIOS_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [92:0] nios_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // NIOS_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> NIOS_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [92:0] nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [92:0] ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_001:sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [92:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_002:sink_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // PCU_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // PCU_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // PCU_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [92:0] pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // PCU_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_003:sink_ready -> PCU_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [92:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // SYSID_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_004:sink_ready -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [92:0] receive_req_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         receive_req_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_005:sink_ready -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [92:0] receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_006:sink_ready -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         req_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // REQ_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         req_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // REQ_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         req_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // REQ_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [92:0] req_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // REQ_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         req_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_007:sink_ready -> REQ_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // ACK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // ACK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // ACK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [92:0] ack_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // ACK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         ack_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> ACK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                              // rst_controller:reset_out -> [NIOS:reset_n, NIOS_data_master_translator:reset, NIOS_data_master_translator_avalon_universal_master_0_agent:reset, NIOS_instruction_master_translator:reset, NIOS_instruction_master_translator_avalon_universal_master_0_agent:reset, NIOS_jtag_debug_module_translator:reset, NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, irq_mapper:reset, rsp_xbar_demux:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset]
	wire         rst_controller_001_reset_out_reset;                                                          // rst_controller_001:reset_out -> [ACK:reset_n, ACK_s1_translator:reset, ACK_s1_translator_avalon_universal_slave_0_agent:reset, ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG:rst_n, JTAG_avalon_jtag_slave_translator:reset, JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PCU:reset_n, PCU_control_slave_translator:reset, PCU_control_slave_translator_avalon_universal_slave_0_agent:reset, PCU_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RAM:reset, RAM_s1_translator:reset, RAM_s1_translator_avalon_universal_slave_0_agent:reset, RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RECEIVE_ACK:reset_n, RECEIVE_ACK_s1_translator:reset, RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:reset, RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RECEIVE_REQ:reset_n, RECEIVE_REQ_s1_translator:reset, RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:reset, RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, REQ:reset_n, REQ_s1_translator:reset, REQ_s1_translator_avalon_universal_slave_0_agent:reset, REQ_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SYSID:reset_n, SYSID_control_slave_translator:reset, SYSID_control_slave_translator_avalon_universal_slave_0_agent:reset, SYSID_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_001:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset]
	wire         nios_jtag_debug_module_reset_reset;                                                          // NIOS:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                             // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                   // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                           // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src0_data;                                                                    // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [8:0] cmd_xbar_demux_src0_channel;                                                                 // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                   // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                             // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                   // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                           // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src1_data;                                                                    // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [8:0] cmd_xbar_demux_src1_channel;                                                                 // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                   // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                         // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                               // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                       // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src0_data;                                                                // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src0_channel;                                                             // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                               // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                         // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                               // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                       // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src1_data;                                                                // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src1_channel;                                                             // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                               // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                         // cmd_xbar_demux_001:src2_endofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                               // cmd_xbar_demux_001:src2_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                       // cmd_xbar_demux_001:src2_startofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src2_data;                                                                // cmd_xbar_demux_001:src2_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src2_channel;                                                             // cmd_xbar_demux_001:src2_channel -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                         // cmd_xbar_demux_001:src3_endofpacket -> PCU_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                               // cmd_xbar_demux_001:src3_valid -> PCU_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                       // cmd_xbar_demux_001:src3_startofpacket -> PCU_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src3_data;                                                                // cmd_xbar_demux_001:src3_data -> PCU_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src3_channel;                                                             // cmd_xbar_demux_001:src3_channel -> PCU_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                         // cmd_xbar_demux_001:src4_endofpacket -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                               // cmd_xbar_demux_001:src4_valid -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                       // cmd_xbar_demux_001:src4_startofpacket -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src4_data;                                                                // cmd_xbar_demux_001:src4_data -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src4_channel;                                                             // cmd_xbar_demux_001:src4_channel -> SYSID_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                         // cmd_xbar_demux_001:src5_endofpacket -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                               // cmd_xbar_demux_001:src5_valid -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                       // cmd_xbar_demux_001:src5_startofpacket -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src5_data;                                                                // cmd_xbar_demux_001:src5_data -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src5_channel;                                                             // cmd_xbar_demux_001:src5_channel -> RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                         // cmd_xbar_demux_001:src6_endofpacket -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                               // cmd_xbar_demux_001:src6_valid -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                       // cmd_xbar_demux_001:src6_startofpacket -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src6_data;                                                                // cmd_xbar_demux_001:src6_data -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src6_channel;                                                             // cmd_xbar_demux_001:src6_channel -> RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                         // cmd_xbar_demux_001:src7_endofpacket -> REQ_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                               // cmd_xbar_demux_001:src7_valid -> REQ_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                       // cmd_xbar_demux_001:src7_startofpacket -> REQ_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src7_data;                                                                // cmd_xbar_demux_001:src7_data -> REQ_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src7_channel;                                                             // cmd_xbar_demux_001:src7_channel -> REQ_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                         // cmd_xbar_demux_001:src8_endofpacket -> ACK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                               // cmd_xbar_demux_001:src8_valid -> ACK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                       // cmd_xbar_demux_001:src8_startofpacket -> ACK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src8_data;                                                                // cmd_xbar_demux_001:src8_data -> ACK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src8_channel;                                                             // cmd_xbar_demux_001:src8_channel -> ACK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                             // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                   // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                           // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_src0_data;                                                                    // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [8:0] rsp_xbar_demux_src0_channel;                                                                 // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                   // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                             // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                   // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                           // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_src1_data;                                                                    // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [8:0] rsp_xbar_demux_src1_channel;                                                                 // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                   // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                         // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                               // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                       // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_001_src0_data;                                                                // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src0_channel;                                                             // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                               // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                         // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                               // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                       // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_001_src1_data;                                                                // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src1_channel;                                                             // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                               // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                         // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                               // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                       // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [92:0] rsp_xbar_demux_002_src0_data;                                                                // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src0_channel;                                                             // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                               // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                         // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                               // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                       // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [92:0] rsp_xbar_demux_003_src0_data;                                                                // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src0_channel;                                                             // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                               // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                         // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                               // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                       // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [92:0] rsp_xbar_demux_004_src0_data;                                                                // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src0_channel;                                                             // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                               // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                         // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                               // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                       // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [92:0] rsp_xbar_demux_005_src0_data;                                                                // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src0_channel;                                                             // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                               // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                         // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                               // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                       // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [92:0] rsp_xbar_demux_006_src0_data;                                                                // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src0_channel;                                                             // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                               // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                         // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                               // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                       // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [92:0] rsp_xbar_demux_007_src0_data;                                                                // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src0_channel;                                                             // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                               // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                         // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                               // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                       // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [92:0] rsp_xbar_demux_008_src0_data;                                                                // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [8:0] rsp_xbar_demux_008_src0_channel;                                                             // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                               // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         addr_router_src_endofpacket;                                                                 // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                       // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                               // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [92:0] addr_router_src_data;                                                                        // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [8:0] addr_router_src_channel;                                                                     // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                       // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                // rsp_xbar_mux:src_endofpacket -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                      // rsp_xbar_mux:src_valid -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                              // rsp_xbar_mux:src_startofpacket -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] rsp_xbar_mux_src_data;                                                                       // rsp_xbar_mux:src_data -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] rsp_xbar_mux_src_channel;                                                                    // rsp_xbar_mux:src_channel -> NIOS_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                      // NIOS_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                             // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                   // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                           // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [92:0] addr_router_001_src_data;                                                                    // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [8:0] addr_router_001_src_channel;                                                                 // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                   // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                            // rsp_xbar_mux_001:src_endofpacket -> NIOS_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                  // rsp_xbar_mux_001:src_valid -> NIOS_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                          // rsp_xbar_mux_001:src_startofpacket -> NIOS_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] rsp_xbar_mux_001_src_data;                                                                   // rsp_xbar_mux_001:src_data -> NIOS_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] rsp_xbar_mux_001_src_channel;                                                                // rsp_xbar_mux_001:src_channel -> NIOS_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                  // NIOS_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                // cmd_xbar_mux:src_endofpacket -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                      // cmd_xbar_mux:src_valid -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                              // cmd_xbar_mux:src_startofpacket -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_src_data;                                                                       // cmd_xbar_mux:src_data -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_src_channel;                                                                    // cmd_xbar_mux:src_channel -> NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                      // NIOS_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                   // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                         // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                 // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [92:0] id_router_src_data;                                                                          // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [8:0] id_router_src_channel;                                                                       // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                         // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                            // cmd_xbar_mux_001:src_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                  // cmd_xbar_mux_001:src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                          // cmd_xbar_mux_001:src_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_001_src_data;                                                                   // cmd_xbar_mux_001:src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_001_src_channel;                                                                // cmd_xbar_mux_001:src_channel -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                  // RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                               // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                     // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                             // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [92:0] id_router_001_src_data;                                                                      // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [8:0] id_router_001_src_channel;                                                                   // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                     // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_001_src2_ready;                                                               // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire         id_router_002_src_endofpacket;                                                               // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                     // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                             // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [92:0] id_router_002_src_data;                                                                      // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [8:0] id_router_002_src_channel;                                                                   // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                     // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                               // PCU_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                               // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                     // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                             // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [92:0] id_router_003_src_data;                                                                      // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [8:0] id_router_003_src_channel;                                                                   // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                     // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                               // SYSID_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                               // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                     // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                             // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [92:0] id_router_004_src_data;                                                                      // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [8:0] id_router_004_src_channel;                                                                   // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                     // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                               // RECEIVE_REQ_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                               // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                     // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                             // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [92:0] id_router_005_src_data;                                                                      // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [8:0] id_router_005_src_channel;                                                                   // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                     // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                               // RECEIVE_ACK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                               // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                     // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                             // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [92:0] id_router_006_src_data;                                                                      // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [8:0] id_router_006_src_channel;                                                                   // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                     // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                               // REQ_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                               // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                     // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                             // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [92:0] id_router_007_src_data;                                                                      // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [8:0] id_router_007_src_channel;                                                                   // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                     // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                               // ACK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                               // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                     // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                             // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [92:0] id_router_008_src_data;                                                                      // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [8:0] id_router_008_src_channel;                                                                   // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                     // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         irq_mapper_receiver0_irq;                                                                    // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_d_irq_irq;                                                                              // irq_mapper:sender_irq -> NIOS:d_irq

	SoC2_NIOS nios (
		.clk                                   (clk_clk),                                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                   //                   reset_n.reset_n
		.d_address                             (nios_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios_data_master_read),                                             //                          .read
		.d_readdata                            (nios_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios_data_master_write),                                            //                          .write
		.d_writedata                           (nios_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                   // custom_instruction_master.readra
	);

	SoC2_RAM ram (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                // reset1.reset
	);

	SoC2_JTAG jtag (
		.clk            (clk_clk),                                                           //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                               //             reset.reset_n
		.av_chipselect  (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                           //               irq.irq
	);

	SoC2_PCU pcu (
		.clk           (clk_clk),                                                        //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                            //         reset.reset_n
		.address       (pcu_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (pcu_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (pcu_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (pcu_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (pcu_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	SoC2_SYSID sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	SoC2_RECEIVE_REQ receive_req (
		.clk      (clk_clk),                                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address  (receive_req_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (receive_req_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (receive_req_export)                                      // external_connection.export
	);

	SoC2_REQ req (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (req_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~req_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (req_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (req_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (req_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (req_export)                                        // external_connection.export
	);

	SoC2_RECEIVE_REQ receive_ack (
		.clk      (clk_clk),                                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address  (receive_ack_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (receive_ack_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (receive_ack_export)                                      // external_connection.export
	);

	SoC2_REQ ack (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (ack_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ack_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ack_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ack_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ack_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ack_export)                                        // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios_instruction_master_translator (
		.clk                      (clk_clk),                                                                    //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                             //                     reset.reset
		.uav_address              (nios_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios_instruction_master_read),                                               //                          .read
		.av_readdata              (nios_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                       //               (terminated)
		.av_byteenable            (4'b1111),                                                                    //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                       //               (terminated)
		.av_begintransfer         (1'b0),                                                                       //               (terminated)
		.av_chipselect            (1'b0),                                                                       //               (terminated)
		.av_readdatavalid         (),                                                                           //               (terminated)
		.av_write                 (1'b0),                                                                       //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                       //               (terminated)
		.av_lock                  (1'b0),                                                                       //               (terminated)
		.av_debugaccess           (1'b0),                                                                       //               (terminated)
		.uav_clken                (),                                                                           //               (terminated)
		.av_clken                 (1'b1),                                                                       //               (terminated)
		.uav_response             (2'b00),                                                                      //               (terminated)
		.av_response              (),                                                                           //               (terminated)
		.uav_writeresponserequest (),                                                                           //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                       //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                       //               (terminated)
		.av_writeresponsevalid    ()                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios_data_master_translator (
		.clk                      (clk_clk),                                                             //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address              (nios_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios_data_master_read),                                               //                          .read
		.av_readdata              (nios_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios_data_master_write),                                              //                          .write
		.av_writedata             (nios_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                //               (terminated)
		.av_begintransfer         (1'b0),                                                                //               (terminated)
		.av_chipselect            (1'b0),                                                                //               (terminated)
		.av_readdatavalid         (),                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                //               (terminated)
		.uav_clken                (),                                                                    //               (terminated)
		.av_clken                 (1'b1),                                                                //               (terminated)
		.uav_response             (2'b00),                                                               //               (terminated)
		.av_response              (),                                                                    //               (terminated)
		.uav_writeresponserequest (),                                                                    //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                //               (terminated)
		.av_writeresponsevalid    ()                                                                     //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_chipselect            (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (14),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address              (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pcu_control_slave_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pcu_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pcu_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pcu_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pcu_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (pcu_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read                  (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) receive_req_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (receive_req_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (receive_req_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_writedata             (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) receive_ack_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (receive_ack_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (receive_ack_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_writedata             (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) req_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (req_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (req_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (req_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (req_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (req_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (req_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (req_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (req_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (req_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (req_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (req_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (req_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (req_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (req_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (req_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (req_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ack_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (ack_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ack_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ack_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ack_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ack_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ack_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ack_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ack_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ack_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                             //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.av_address              (nios_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                              //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                               //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                            //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                              //          .ready
		.av_response             (),                                                                                    // (terminated)
		.av_writeresponserequest (1'b0),                                                                                // (terminated)
		.av_writeresponsevalid   ()                                                                                     // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                      //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address              (nios_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                   //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                    //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                 //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                             //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                   //          .ready
		.av_response             (),                                                                             // (terminated)
		.av_writeresponserequest (1'b0),                                                                         // (terminated)
		.av_writeresponsevalid   ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                    //                .channel
		.rf_sink_ready           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                //                .channel
		.rf_sink_ready           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                             //                .channel
		.rf_sink_ready           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pcu_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pcu_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                        //                .channel
		.rf_sink_ready           (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pcu_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pcu_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pcu_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) receive_req_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (receive_req_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                     //                .channel
		.rf_sink_ready           (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (receive_req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (receive_req_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (receive_req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) receive_ack_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (receive_ack_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                     //                .channel
		.rf_sink_ready           (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (receive_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (receive_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (receive_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) req_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (req_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (req_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (req_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (req_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (req_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (req_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (req_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (req_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (req_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (req_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (req_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (req_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (req_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (req_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (req_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (req_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                             //                .channel
		.rf_sink_ready           (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (req_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (req_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (req_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (req_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (req_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (req_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (req_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (req_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (req_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (req_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (req_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (req_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ack_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (ack_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ack_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ack_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ack_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ack_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ack_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ack_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                             //                .channel
		.rf_sink_ready           (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	SoC2_addr_router addr_router (
		.sink_ready         (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_src_valid),                                                               //          .valid
		.src_data           (addr_router_src_data),                                                                //          .data
		.src_channel        (addr_router_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                          //          .endofpacket
	);

	SoC2_addr_router_001 addr_router_001 (
		.sink_ready         (nios_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                    //          .valid
		.src_data           (addr_router_001_src_data),                                                     //          .data
		.src_channel        (addr_router_001_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                               //          .endofpacket
	);

	SoC2_id_router id_router (
		.sink_ready         (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                               //       src.ready
		.src_valid          (id_router_src_valid),                                                               //          .valid
		.src_data           (id_router_src_data),                                                                //          .data
		.src_channel        (id_router_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                          //          .endofpacket
	);

	SoC2_id_router id_router_001 (
		.sink_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                           //          .valid
		.src_data           (id_router_001_src_data),                                            //          .data
		.src_channel        (id_router_001_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                      //          .endofpacket
	);

	SoC2_id_router_002 id_router_002 (
		.sink_ready         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                                           //          .valid
		.src_data           (id_router_002_src_data),                                                            //          .data
		.src_channel        (id_router_002_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                      //          .endofpacket
	);

	SoC2_id_router_002 id_router_003 (
		.sink_ready         (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcu_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                      //       src.ready
		.src_valid          (id_router_003_src_valid),                                                      //          .valid
		.src_data           (id_router_003_src_data),                                                       //          .data
		.src_channel        (id_router_003_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                 //          .endofpacket
	);

	SoC2_id_router_002 id_router_004 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                        //       src.ready
		.src_valid          (id_router_004_src_valid),                                                        //          .valid
		.src_data           (id_router_004_src_data),                                                         //          .data
		.src_channel        (id_router_004_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                   //          .endofpacket
	);

	SoC2_id_router_002 id_router_005 (
		.sink_ready         (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (receive_req_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                   //       src.ready
		.src_valid          (id_router_005_src_valid),                                                   //          .valid
		.src_data           (id_router_005_src_data),                                                    //          .data
		.src_channel        (id_router_005_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                              //          .endofpacket
	);

	SoC2_id_router_002 id_router_006 (
		.sink_ready         (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (receive_ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                   //       src.ready
		.src_valid          (id_router_006_src_valid),                                                   //          .valid
		.src_data           (id_router_006_src_data),                                                    //          .data
		.src_channel        (id_router_006_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                              //          .endofpacket
	);

	SoC2_id_router_002 id_router_007 (
		.sink_ready         (req_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (req_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (req_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (req_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (req_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                           //       src.ready
		.src_valid          (id_router_007_src_valid),                                           //          .valid
		.src_data           (id_router_007_src_data),                                            //          .data
		.src_channel        (id_router_007_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                      //          .endofpacket
	);

	SoC2_id_router_002 id_router_008 (
		.sink_ready         (ack_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ack_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ack_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                           //       src.ready
		.src_valid          (id_router_008_src_valid),                                           //          .valid
		.src_data           (id_router_008_src_data),                                            //          .data
		.src_channel        (id_router_008_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                      //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (nios_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	SoC2_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	SoC2_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),         //      src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	SoC2_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC2_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SoC2_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	SoC2_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SoC2_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	SoC2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_d_irq_irq)                  //    sender.irq
	);

endmodule
